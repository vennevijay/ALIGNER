`define CFS_ALGN_TEST_ALGN_DATA_WIDTH 32